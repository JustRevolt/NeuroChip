`define VIVADO_PRJ_USE
`define DEBUG